module fd_reg(pc_in, ir_in, pc_out, ir_out, clk, clear);

	input [31:0] pc_in, ir_in;
	input clk, clear;
	output [31:0] pc_out, ir_out;
	
	flip_floppity_flop pc_0(pc_out[0], pc_in[0], clk, clear);
	flip_floppity_flop pc_1(pc_out[1], pc_in[1], clk, clear);
	flip_floppity_flop pc_2(pc_out[2], pc_in[2], clk, clear);
	flip_floppity_flop pc_3(pc_out[3], pc_in[3], clk, clear);
	flip_floppity_flop pc_4(pc_out[4], pc_in[4], clk, clear);
	flip_floppity_flop pc_5(pc_out[5], pc_in[5], clk, clear);
	flip_floppity_flop pc_6(pc_out[6], pc_in[6], clk, clear);
	flip_floppity_flop pc_7(pc_out[7], pc_in[7], clk, clear);
	flip_floppity_flop pc_8(pc_out[8], pc_in[8], clk, clear);
	flip_floppity_flop pc_9(pc_out[9], pc_in[9], clk, clear);
	flip_floppity_flop pc_10(pc_out[10], pc_in[10], clk, clear);
	flip_floppity_flop pc_11(pc_out[11], pc_in[11], clk, clear);
	flip_floppity_flop pc_12(pc_out[12], pc_in[12], clk, clear);
	flip_floppity_flop pc_13(pc_out[13], pc_in[13], clk, clear);
	flip_floppity_flop pc_14(pc_out[14], pc_in[14], clk, clear);
	flip_floppity_flop pc_15(pc_out[15], pc_in[15], clk, clear);
	flip_floppity_flop pc_16(pc_out[16], pc_in[16], clk, clear);
	flip_floppity_flop pc_17(pc_out[17], pc_in[17], clk, clear);
	flip_floppity_flop pc_18(pc_out[18], pc_in[18], clk, clear);
	flip_floppity_flop pc_19(pc_out[19], pc_in[19], clk, clear);
	flip_floppity_flop pc_20(pc_out[20], pc_in[20], clk, clear);
	flip_floppity_flop pc_21(pc_out[21], pc_in[21], clk, clear);
	flip_floppity_flop pc_22(pc_out[22], pc_in[22], clk, clear);
	flip_floppity_flop pc_23(pc_out[23], pc_in[23], clk, clear);
	flip_floppity_flop pc_24(pc_out[24], pc_in[24], clk, clear);
	flip_floppity_flop pc_25(pc_out[25], pc_in[25], clk, clear);
	flip_floppity_flop pc_26(pc_out[26], pc_in[26], clk, clear);
	flip_floppity_flop pc_27(pc_out[27], pc_in[27], clk, clear);
	flip_floppity_flop pc_28(pc_out[28], pc_in[28], clk, clear);
	flip_floppity_flop pc_29(pc_out[29], pc_in[29], clk, clear);
	flip_floppity_flop pc_30(pc_out[30], pc_in[30], clk, clear);
	flip_floppity_flop pc_31(pc_out[31], pc_in[31], clk, clear);
	
	flip_floppity_flop ir_0(ir_out[0], ir_in[0], clk, clear);
	flip_floppity_flop ir_1(ir_out[1], ir_in[1], clk, clear);
	flip_floppity_flop ir_2(ir_out[2], ir_in[2], clk, clear);
	flip_floppity_flop ir_3(ir_out[3], ir_in[3], clk, clear);
	flip_floppity_flop ir_4(ir_out[4], ir_in[4], clk, clear);
	flip_floppity_flop ir_5(ir_out[5], ir_in[5], clk, clear);
	flip_floppity_flop ir_6(ir_out[6], ir_in[6], clk, clear);
	flip_floppity_flop ir_7(ir_out[7], ir_in[7], clk, clear);
	flip_floppity_flop ir_8(ir_out[8], ir_in[8], clk, clear);
	flip_floppity_flop ir_9(ir_out[9], ir_in[9], clk, clear);
	flip_floppity_flop ir_10(ir_out[10], ir_in[10], clk, clear);
	flip_floppity_flop ir_11(ir_out[11], ir_in[11], clk, clear);
	flip_floppity_flop ir_12(ir_out[12], ir_in[12], clk, clear);
	flip_floppity_flop ir_13(ir_out[13], ir_in[13], clk, clear);
	flip_floppity_flop ir_14(ir_out[14], ir_in[14], clk, clear);
	flip_floppity_flop ir_15(ir_out[15], ir_in[15], clk, clear);
	flip_floppity_flop ir_16(ir_out[16], ir_in[16], clk, clear);
	flip_floppity_flop ir_17(ir_out[17], ir_in[17], clk, clear);
	flip_floppity_flop ir_18(ir_out[18], ir_in[18], clk, clear);
	flip_floppity_flop ir_19(ir_out[19], ir_in[19], clk, clear);
	flip_floppity_flop ir_20(ir_out[20], ir_in[20], clk, clear);
	flip_floppity_flop ir_21(ir_out[21], ir_in[21], clk, clear);
	flip_floppity_flop ir_22(ir_out[22], ir_in[22], clk, clear);
	flip_floppity_flop ir_23(ir_out[23], ir_in[23], clk, clear);
	flip_floppity_flop ir_24(ir_out[24], ir_in[24], clk, clear);
	flip_floppity_flop ir_25(ir_out[25], ir_in[25], clk, clear);
	flip_floppity_flop ir_26(ir_out[26], ir_in[26], clk, clear);
	flip_floppity_flop ir_27(ir_out[27], ir_in[27], clk, clear);
	flip_floppity_flop ir_28(ir_out[28], ir_in[28], clk, clear);
	flip_floppity_flop ir_29(ir_out[29], ir_in[29], clk, clear);
	flip_floppity_flop ir_30(ir_out[30], ir_in[30], clk, clear);
	flip_floppity_flop ir_31(ir_out[31], ir_in[31], clk, clear);
	
endmodule
