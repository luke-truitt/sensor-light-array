module test_loop(out, in);

	input[31:0]