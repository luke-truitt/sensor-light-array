module and_32(out, in1, in2);
	
	input [31:0] in1, in2;
	output [31:0] out;
	
	and and1(out, in1, in2);
	
endmodule;
