module reg_64(out, in, clk, clear);

input [63:0] in;
	input clk, clear;
	output [63:0] out;
	
	flip_floppity_flop dff_0(out[0], in[0], clk, clear);
	flip_floppity_flop dff_1(out[1], in[1], clk, clear);
	flip_floppity_flop dff_2(out[2], in[2], clk, clear);
	flip_floppity_flop dff_3(out[3], in[3], clk, clear);
	flip_floppity_flop dff_4(out[4], in[4], clk, clear);
	flip_floppity_flop dff_5(out[5], in[5], clk, clear);
	flip_floppity_flop dff_6(out[6], in[6], clk, clear);
	flip_floppity_flop dff_7(out[7], in[7], clk, clear);
	flip_floppity_flop dff_8(out[8], in[8], clk, clear);
	flip_floppity_flop dff_9(out[9], in[9], clk, clear);
	flip_floppity_flop dff_10(out[10], in[10], clk, clear);
	flip_floppity_flop dff_11(out[11], in[11], clk, clear);
	flip_floppity_flop dff_12(out[12], in[12], clk, clear);
	flip_floppity_flop dff_13(out[13], in[13], clk, clear);
	flip_floppity_flop dff_14(out[14], in[14], clk, clear);
	flip_floppity_flop dff_15(out[15], in[15], clk, clear);
	flip_floppity_flop dff_16(out[16], in[16], clk, clear);
	flip_floppity_flop dff_17(out[17], in[17], clk, clear);
	flip_floppity_flop dff_18(out[18], in[18], clk, clear);
	flip_floppity_flop dff_19(out[19], in[19], clk, clear);
	flip_floppity_flop dff_20(out[20], in[20], clk, clear);
	flip_floppity_flop dff_21(out[21], in[21], clk, clear);
	flip_floppity_flop dff_22(out[22], in[22], clk, clear);
	flip_floppity_flop dff_23(out[23], in[23], clk, clear);
	flip_floppity_flop dff_24(out[24], in[24], clk, clear);
	flip_floppity_flop dff_25(out[25], in[25], clk, clear);
	flip_floppity_flop dff_26(out[26], in[26], clk, clear);
	flip_floppity_flop dff_27(out[27], in[27], clk, clear);
	flip_floppity_flop dff_28(out[28], in[28], clk, clear);
	flip_floppity_flop dff_29(out[29], in[29], clk, clear);
	flip_floppity_flop dff_30(out[30], in[30], clk, clear);
	flip_floppity_flop dff_31(out[31], in[31], clk, clear);
	flip_floppity_flop dff_32(out[32], in[32], clk, clear);
	flip_floppity_flop dff_33(out[33], in[33], clk, clear);
	flip_floppity_flop dff_34(out[34], in[34], clk, clear);
	flip_floppity_flop dff_35(out[35], in[35], clk, clear);
	flip_floppity_flop dff_36(out[36], in[36], clk, clear);
	flip_floppity_flop dff_37(out[37], in[37], clk, clear);
	flip_floppity_flop dff_38(out[38], in[38], clk, clear);
	flip_floppity_flop dff_39(out[39], in[39], clk, clear);
	flip_floppity_flop dff_40(out[40], in[40], clk, clear);
	flip_floppity_flop dff_41(out[41], in[41], clk, clear);
	flip_floppity_flop dff_42(out[42], in[42], clk, clear);
	flip_floppity_flop dff_43(out[43], in[43], clk, clear);
	flip_floppity_flop dff_44(out[44], in[44], clk, clear);
	flip_floppity_flop dff_45(out[45], in[45], clk, clear);
	flip_floppity_flop dff_46(out[46], in[46], clk, clear);
	flip_floppity_flop dff_47(out[47], in[47], clk, clear);
	flip_floppity_flop dff_48(out[48], in[48], clk, clear);
	flip_floppity_flop dff_49(out[49], in[49], clk, clear);
	flip_floppity_flop dff_50(out[50], in[50], clk, clear);
	flip_floppity_flop dff_51(out[51], in[51], clk, clear);
	flip_floppity_flop dff_52(out[52], in[52], clk, clear);
	flip_floppity_flop dff_53(out[53], in[53], clk, clear);
	flip_floppity_flop dff_54(out[54], in[54], clk, clear);
	flip_floppity_flop dff_55(out[55], in[55], clk, clear);
	flip_floppity_flop dff_56(out[56], in[56], clk, clear);
	flip_floppity_flop dff_57(out[57], in[57], clk, clear);
	flip_floppity_flop dff_58(out[58], in[58], clk, clear);
	flip_floppity_flop dff_59(out[59], in[59], clk, clear);
	flip_floppity_flop dff_60(out[60], in[60], clk, clear);
	flip_floppity_flop dff_61(out[61], in[61], clk, clear);
	flip_floppity_flop dff_62(out[62], in[62], clk, clear);
	flip_floppity_flop dff_63(out[63], in[63], clk, clear);
	
endmodule
